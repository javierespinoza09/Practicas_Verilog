module RegistroControl2 (
    input CLK, EN, RESET,
    input [31:0] GENERADOR_DATOS, REGISTRO_DATOS,
    output FLAG, NEW,    
    
    //VARIABLES SOLAMENTE PARA LA COMPORBACION DE LA SIMULACION 
    //DEBEN IR COMENTADAS
    output [11:0] COMPARADOR_DATOS, //ESTA ENTRADA BORRARLA, SOLAMENTE SE NECESITA, PARA REALIZAR LAS DIVERSAS SIMULACIONES DE COMPARACION.
    output [11:0] UMBRAL //ESTA ENTRADA BORRARLA, SOLAMENTE SE NECESITA, PARA REALIZAR LAS DIVERSAS SIMULACIONES DE COMPARACION.
    );
    
    reg [31:0] REGISTRO_CONTROL;
    reg [11:0] COMPARADOR_REGISTRO_DATOS;
    reg [11:0] UMBRAL_GENERADOR_DATOS;
    
    always @(posedge CLK)begin
        if(EN == 1) begin
            if(RESET == 1) REGISTRO_CONTROL <= 32'b0; //RESET ACTIVADO EN ALTO
            else begin
            REGISTRO_CONTROL[15:8] <= GENERADOR_DATOS[15:8]; //SE ASIGNA EL VALOR DEL UMBRAL
            UMBRAL_GENERADOR_DATOS <= REGISTRO_CONTROL[15:8] << 4; //SE REALIZA EL CORRIMIENTO DE 4 BITS           
            COMPARADOR_REGISTRO_DATOS <= REGISTRO_DATOS[11:0]; //SE ASIGNA EL VALOR A COMPARAR DEL ADC
            
            //COLOCA EL FLAG
            if(COMPARADOR_REGISTRO_DATOS > UMBRAL_GENERADOR_DATOS) REGISTRO_CONTROL[1] = 1;
            else if(COMPARADOR_REGISTRO_DATOS < UMBRAL_GENERADOR_DATOS) REGISTRO_CONTROL[1] = 0;    
            
            //COLOCA EL NEW
            if (REGISTRO_CONTROL[0] == 1) REGISTRO_CONTROL[0] <= 0; //SE RESTABLECE EL NEW
            else REGISTRO_CONTROL[0] <= GENERADOR_DATOS[0]; //SE ESTABLECE EL NEW
            
            end 
        end
    end
    
    assign FLAG = REGISTRO_CONTROL[1];
    assign NEW = REGISTRO_CONTROL[0];  
    
    //VARIABLES SOLAMENTE PARA LA COMPORBACION DE LA SIMULACION 
    //DEBEN IR COMENTADAS
    assign COMPARADOR_DATOS = COMPARADOR_REGISTRO_DATOS; // ESTA ENTRADA BORRARLA, SOLAMENTE SE NECESITA, PARA REALIZAR LAS DIVERSAS SIMULACIONES DE COMPARACION.
    assign UMBRAL = UMBRAL_GENERADOR_DATOS; // ESTA ENTRADA BORRARLA, SOLAMENTE SE NECESITA, PARA REALIZAR LAS DIVERSAS SIMULACIONES DE COMPARACION.      
       
endmodule