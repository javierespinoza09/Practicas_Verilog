module ak7();
endmodule
