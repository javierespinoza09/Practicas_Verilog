module 
endmodule
