// Code your design here
module f (input [3:0] a, output reg [3:0] b);
  assign b = a+1;
  
endmodule 